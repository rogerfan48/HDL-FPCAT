module game_engine(
    
);

endmodule